magic
tech sky130A
magscale 1 2
timestamp 1729313229
<< viali >>
rect 1070 1511 1122 1563
<< metal1 >>
rect -244 2743 1579 2789
rect 972 2369 1018 2371
rect 1110 2369 1156 2604
rect 1533 2372 1579 2743
rect 972 2323 1383 2369
rect 972 2321 1018 2323
rect 1009 2059 1015 2062
rect 884 2013 1015 2059
rect 1009 2010 1015 2013
rect 1067 2010 1073 2062
rect 1084 1691 1442 1720
rect 230 1453 276 1620
rect 1084 1569 1113 1691
rect 1430 1651 1432 1660
rect 1185 1622 1434 1651
rect 1058 1563 1134 1569
rect 1058 1511 1070 1563
rect 1122 1511 1134 1563
rect 1058 1505 1134 1511
rect 1185 1477 1215 1622
rect 1430 1614 1432 1622
rect 230 1407 539 1453
rect 1060 1425 1070 1477
rect 1122 1425 1215 1477
rect -522 1354 15 1400
rect -43 1151 15 1354
rect 493 1240 539 1407
rect -393 826 -177 872
rect -207 137 -177 826
rect -207 91 -31 137
<< via1 >>
rect 1015 2010 1067 2062
rect 1070 1425 1122 1477
<< metal2 >>
rect 1017 2068 1063 2604
rect 1015 2062 1067 2068
rect 1067 2013 1335 2059
rect 1015 2004 1067 2010
rect 1442 1599 1510 1675
rect 1070 1477 1122 1487
rect -156 1459 -147 1461
rect -391 1403 -147 1459
rect -156 1401 -147 1403
rect -87 1401 -78 1461
rect 1070 1415 1122 1425
rect 375 1067 427 1398
<< via2 >>
rect -147 1401 -87 1461
<< metal3 >>
rect 1517 1604 1520 1670
rect -152 1461 -82 1466
rect -152 1401 -147 1461
rect -87 1401 1593 1461
rect -152 1396 -82 1401
use nmos34  nmos34_0
timestamp 1729220844
transform 1 0 115 0 -1 1167
box -292 -79 984 1161
use nmos89  nmos89_0
timestamp 1729243167
transform 1 0 -84 0 -1 2023
box -93 -433 1201 409
use pmos67  pmos67_0
timestamp 1729238107
transform 1 0 1344 0 1 1755
box -197 -1743 621 693
use pmoscs  pmoscs_0
timestamp 1729159655
transform 1 0 -1021 0 1 815
box -189 -803 814 2080
<< labels >>
flabel metal1 518 2764 518 2764 0 FreeSans 1600 0 0 0 VDD
port 0 nsew
flabel viali 1092 1536 1092 1536 0 FreeSans 1600 0 0 0 VIP
port 1 nsew
flabel via1 1084 1468 1084 1468 0 FreeSans 1600 0 0 0 VIN
port 2 nsew
flabel metal1 518 1354 518 1354 0 FreeSans 1600 0 0 0 GND
port 3 nsew
flabel metal2 400 1364 400 1364 0 FreeSans 1600 0 0 0 RS
port 4 nsew
flabel metal1 1134 2586 1134 2586 0 FreeSans 1600 0 0 0 OUT
port 5 nsew
<< end >>
