magic
tech sky130A
magscale 1 2
timestamp 1729223874
<< psubdiff >>
rect -293 625 -233 659
rect 931 625 991 659
rect -293 599 -259 625
rect 957 599 991 625
rect -293 -547 -259 -521
rect 957 -547 991 -521
rect -293 -581 -233 -547
rect 931 -581 991 -547
<< psubdiffcont >>
rect -233 625 931 659
rect -293 -521 -259 599
rect 957 -521 991 599
rect -233 -581 931 -547
<< poly >>
rect 253 515 449 576
rect 250 4 451 64
rect 252 -510 448 -449
<< locali >>
rect -293 625 -233 659
rect 931 625 991 659
rect -293 599 -259 625
rect -293 -547 -259 -521
rect 957 599 991 625
rect 957 -547 991 -521
rect -293 -581 -233 -547
rect 931 -581 991 -547
<< viali >>
rect 270 625 304 659
rect 401 -581 435 -547
<< metal1 >>
rect 258 659 316 665
rect 258 625 270 659
rect 304 625 316 659
rect 258 619 316 625
rect -192 470 -158 566
rect -104 477 -70 566
rect -104 470 17 477
rect 270 471 304 619
rect 769 476 803 566
rect 857 479 891 566
rect -78 106 17 470
rect -78 100 46 106
rect 12 56 46 100
rect 12 10 96 56
rect 270 50 304 114
rect 378 101 388 476
rect 440 101 450 476
rect 669 244 803 476
rect 633 153 643 244
rect 705 153 803 244
rect 669 99 803 153
rect 860 470 891 479
rect 860 99 867 470
rect 269 16 430 50
rect -75 -34 18 -33
rect 270 -34 304 -33
rect -75 -404 2 -34
rect -191 -500 -157 -404
rect -103 -410 2 -404
rect 54 -410 64 -34
rect 250 -410 260 -34
rect 312 -410 322 -34
rect 395 -38 430 16
rect 604 10 688 56
rect 654 -33 688 10
rect 654 -40 774 -33
rect 681 -404 774 -40
rect -103 -500 -69 -410
rect 396 -541 430 -404
rect 681 -410 802 -404
rect 768 -500 802 -410
rect 856 -500 890 -404
rect 389 -547 447 -541
rect 389 -581 401 -547
rect 435 -581 447 -547
rect 389 -587 447 -581
<< via1 >>
rect 388 101 440 476
rect 643 153 705 244
rect 2 -410 54 -34
rect 260 -410 312 -34
<< metal2 >>
rect 388 476 440 486
rect 646 476 702 486
rect 643 244 646 254
rect 702 244 705 254
rect 643 143 646 153
rect 388 52 440 101
rect 702 143 705 153
rect 646 91 702 101
rect 259 16 440 52
rect 0 -34 56 -24
rect 0 -420 56 -410
rect 260 -34 312 16
rect 388 15 440 16
rect 260 -420 312 -410
<< via2 >>
rect 646 244 702 476
rect 646 153 702 244
rect 646 101 702 153
rect 0 -410 2 -34
rect 2 -410 54 -34
rect 54 -410 56 -34
<< metal3 >>
rect 636 476 712 481
rect 636 101 646 476
rect 702 101 712 476
rect 636 64 712 101
rect -10 2 712 64
rect -10 -34 66 2
rect 636 1 712 2
rect -10 -410 0 -34
rect 56 -410 66 -34
rect -10 -415 66 -410
use sky130_fd_pr__nfet_01v8_7QRB7N  sky130_fd_pr__nfet_01v8_7QRB7N_0
timestamp 1729218371
transform 1 0 158 0 1 288
box -158 -288 158 288
use sky130_fd_pr__nfet_01v8_46AAJJ  sky130_fd_pr__nfet_01v8_46AAJJ_0
timestamp 1729218371
transform 1 0 158 0 1 -222
box -158 -288 158 288
use sky130_fd_pr__nfet_01v8_46AAJJ  sky130_fd_pr__nfet_01v8_46AAJJ_1
timestamp 1729218371
transform 1 0 542 0 1 -222
box -158 -288 158 288
use sky130_fd_pr__nfet_01v8_46AAJJ  sky130_fd_pr__nfet_01v8_46AAJJ_2
timestamp 1729218371
transform 1 0 542 0 1 288
box -158 -288 158 288
use sky130_fd_pr__nfet_01v8_TCR5KT  sky130_fd_pr__nfet_01v8_TCR5KT_0
timestamp 1729217068
transform -1 0 829 0 -1 -253
box -73 -257 73 257
use sky130_fd_pr__nfet_01v8_TCR5KT  sky130_fd_pr__nfet_01v8_TCR5KT_1
timestamp 1729217068
transform 1 0 -131 0 1 319
box -73 -257 73 257
use sky130_fd_pr__nfet_01v8_TCR5KT  sky130_fd_pr__nfet_01v8_TCR5KT_2
timestamp 1729217068
transform 1 0 830 0 1 319
box -73 -257 73 257
use sky130_fd_pr__nfet_01v8_TCR5KT  sky130_fd_pr__nfet_01v8_TCR5KT_3
timestamp 1729217068
transform -1 0 -130 0 -1 -253
box -73 -257 73 257
<< labels >>
flabel metal1 19 76 21 77 0 FreeSans 800 0 0 0 D1
port 0 nsew
flabel metal2 274 -9 276 -9 0 FreeSans 800 0 0 0 RS
port 1 nsew
flabel metal3 690 68 704 70 0 FreeSans 800 0 0 0 D4
port 2 nsew
flabel metal1 407 -528 407 -528 0 FreeSans 800 0 0 0 GND
port 3 nsew
<< end >>
