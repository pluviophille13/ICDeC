magic
tech sky130A
magscale 1 2
timestamp 1729222752
<< nmos >>
rect -200 -100 200 100
<< ndiff >>
rect -258 88 -200 100
rect -258 -88 -246 88
rect -212 -88 -200 88
rect -258 -100 -200 -88
rect 200 88 258 100
rect 200 -88 212 88
rect 246 -88 258 88
rect 200 -100 258 -88
<< ndiffc >>
rect -246 -88 -212 88
rect 212 -88 246 88
<< poly >>
rect -200 172 200 188
rect -200 138 -184 172
rect 184 138 200 172
rect -200 100 200 138
rect -200 -138 200 -100
rect -200 -172 -184 -138
rect 184 -172 200 -138
rect -200 -188 200 -172
<< polycont >>
rect -184 138 184 172
rect -184 -172 184 -138
<< locali >>
rect -200 138 -184 172
rect 184 138 200 172
rect -246 88 -212 104
rect -246 -104 -212 -88
rect 212 88 246 104
rect 212 -104 246 -88
rect -200 -172 -184 -138
rect 184 -172 200 -138
<< viali >>
rect -129 138 129 172
rect -246 -88 -212 88
rect 212 -88 246 88
rect -129 -172 129 -138
<< metal1 >>
rect -141 172 141 178
rect -141 138 -129 172
rect 129 138 141 172
rect -141 132 141 138
rect -252 88 -206 100
rect -252 -88 -246 88
rect -212 -88 -206 88
rect -252 -100 -206 -88
rect 206 88 252 100
rect 206 -88 212 88
rect 246 -88 252 88
rect 206 -100 252 -88
rect -141 -138 141 -132
rect -141 -172 -129 -138
rect 129 -172 141 -138
rect -141 -178 141 -172
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1 l 2 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 1 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 70 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
