magic
tech sky130A
timestamp 1729225432
<< nmos >>
rect -25 -40 25 40
<< ndiff >>
rect -54 34 -25 40
rect -54 -34 -48 34
rect -31 -34 -25 34
rect -54 -40 -25 -34
rect 25 34 54 40
rect 25 -34 31 34
rect 48 -34 54 34
rect 25 -40 54 -34
<< ndiffc >>
rect -48 -34 -31 34
rect 31 -34 48 34
<< poly >>
rect -25 76 25 84
rect -25 59 -17 76
rect 17 59 25 76
rect -25 40 25 59
rect -25 -59 25 -40
rect -25 -76 -17 -59
rect 17 -76 25 -59
rect -25 -84 25 -76
<< polycont >>
rect -17 59 17 76
rect -17 -76 17 -59
<< locali >>
rect -25 59 -17 76
rect 17 59 25 76
rect -48 34 -31 42
rect -48 -42 -31 -34
rect 31 34 48 42
rect 31 -42 48 -34
rect -25 -76 -17 -59
rect 17 -76 25 -59
<< viali >>
rect -17 59 17 76
rect -48 -34 -31 34
rect 31 -34 48 34
rect -17 -76 17 -59
<< metal1 >>
rect -23 76 23 79
rect -23 59 -17 76
rect 17 59 23 76
rect -23 56 23 59
rect -51 34 -28 40
rect -51 -34 -48 34
rect -31 -34 -28 34
rect -51 -40 -28 -34
rect 28 34 51 40
rect 28 -34 31 34
rect 48 -34 51 34
rect 28 -40 51 -34
rect -23 -59 23 -56
rect -23 -76 -17 -59
rect 17 -76 23 -59
rect -23 -79 23 -76
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.8 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 1 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
