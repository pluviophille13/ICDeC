magic
tech sky130A
magscale 1 2
timestamp 1729242611
<< psubdiff >>
rect -146 -338 -86 -304
rect 1076 -338 1136 -304
rect -146 -364 -112 -338
rect 1102 -364 1136 -338
rect -146 -1087 -112 -1061
rect 1102 -1087 1136 -1061
rect -146 -1121 -86 -1087
rect 1076 -1121 1136 -1087
<< psubdiffcont >>
rect -86 -338 1076 -304
rect -146 -1061 -112 -364
rect 1102 -1061 1136 -364
rect -86 -1121 1076 -1087
<< poly >>
rect -62 -385 30 -369
rect -62 -419 -46 -385
rect -12 -419 30 -385
rect -62 -435 30 -419
rect 960 -385 1052 -369
rect 960 -419 1002 -385
rect 1036 -419 1052 -385
rect 960 -435 1052 -419
rect 0 -989 30 -980
rect -62 -1005 30 -989
rect -62 -1039 -46 -1005
rect -12 -1039 30 -1005
rect -62 -1055 30 -1039
rect 960 -989 990 -987
rect 960 -1005 1052 -989
rect 960 -1039 1002 -1005
rect 1036 -1039 1052 -1005
rect 960 -1055 1052 -1039
<< polycont >>
rect -46 -419 -12 -385
rect 1002 -419 1036 -385
rect -46 -1039 -12 -1005
rect 1002 -1039 1036 -1005
<< locali >>
rect -146 -338 -86 -304
rect 1076 -338 1136 -304
rect -146 -364 -112 -338
rect 1102 -364 1136 -338
rect -62 -419 -46 -385
rect -12 -419 4 -385
rect 986 -419 1002 -385
rect 1036 -419 1052 -385
rect -46 -465 -12 -419
rect 1002 -464 1036 -419
rect -46 -1005 -12 -960
rect 1001 -1005 1036 -962
rect -62 -1039 -46 -1005
rect -12 -1039 4 -1005
rect 986 -1039 1002 -1005
rect 1036 -1039 1052 -1005
rect -146 -1087 -112 -1061
rect 1102 -1087 1136 -1061
rect -146 -1121 -86 -1087
rect 1076 -1121 1136 -1087
<< viali >>
rect 260 -338 294 -304
rect 696 -338 730 -304
rect -46 -419 -12 -385
rect 1002 -419 1036 -385
rect -46 -1039 -12 -1005
rect 1002 -1039 1036 -1005
rect 260 -1121 294 -1087
rect 696 -1121 730 -1088
rect 696 -1122 730 -1121
<< metal1 >>
rect 248 -304 306 -298
rect 248 -338 260 -304
rect 294 -338 306 -304
rect 248 -344 306 -338
rect 684 -304 742 -298
rect 684 -338 696 -304
rect 730 -338 742 -304
rect 684 -344 742 -338
rect -58 -385 0 -379
rect -58 -419 -46 -385
rect -12 -419 0 -385
rect -58 -425 0 -419
rect -46 -465 -12 -425
rect 257 -466 296 -344
rect 693 -467 732 -344
rect 990 -385 1048 -379
rect 990 -419 1002 -385
rect 1036 -419 1048 -385
rect 990 -425 1048 -419
rect 1002 -464 1036 -425
rect -44 -645 76 -472
rect -44 -646 77 -645
rect 459 -646 469 -469
rect 521 -646 531 -469
rect 915 -644 1035 -470
rect 42 -689 77 -646
rect 914 -689 949 -647
rect 42 -735 949 -689
rect 477 -779 513 -735
rect 22 -782 32 -779
rect -49 -954 32 -782
rect 84 -954 94 -779
rect -49 -956 71 -954
rect 895 -955 905 -778
rect 957 -781 967 -778
rect 957 -955 1033 -781
rect -46 -999 -12 -960
rect -58 -1005 0 -999
rect -58 -1039 -46 -1005
rect -12 -1039 0 -1005
rect -58 -1046 0 -1039
rect 258 -1081 297 -959
rect 248 -1087 306 -1081
rect 693 -1082 732 -958
rect 1001 -999 1036 -962
rect 990 -1005 1048 -999
rect 990 -1039 1002 -1005
rect 1036 -1039 1048 -1005
rect 990 -1045 1048 -1039
rect 248 -1121 260 -1087
rect 294 -1121 306 -1087
rect 248 -1127 306 -1121
rect 684 -1088 742 -1082
rect 684 -1122 696 -1088
rect 730 -1122 742 -1088
rect 684 -1128 742 -1122
<< via1 >>
rect 469 -646 521 -469
rect 32 -954 84 -779
rect 905 -955 957 -778
<< metal2 >>
rect 469 -469 521 -459
rect 469 -688 521 -646
rect 32 -737 958 -688
rect 32 -779 84 -737
rect 32 -964 84 -954
rect 905 -767 958 -737
rect 905 -778 957 -767
rect 905 -965 957 -955
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_0
timestamp 1729225432
transform 1 0 975 0 1 -867
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_1
timestamp 1729225432
transform 1 0 15 0 1 -557
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_2
timestamp 1729225432
transform 1 0 15 0 1 -867
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_3
timestamp 1729225432
transform 1 0 975 0 1 -557
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_YYNGNX  sky130_fd_pr__nfet_01v8_YYNGNX_0
timestamp 1729233197
transform 1 0 495 0 1 -712
box -465 -343 465 343
<< labels >>
flabel metal1 135 -601 197 -535 0 FreeSans 160 0 0 0 M8
flabel metal1 789 -601 851 -535 0 FreeSans 160 0 0 0 M8
flabel metal1 562 -907 624 -841 0 FreeSans 160 0 0 0 M8
flabel metal1 358 -907 420 -841 0 FreeSans 160 0 0 0 M8
flabel metal1 571 -603 633 -537 0 FreeSans 160 0 0 0 M9
flabel metal1 353 -601 415 -535 0 FreeSans 160 0 0 0 M9
flabel metal1 797 -911 859 -845 0 FreeSans 160 0 0 0 M9
flabel metal1 139 -908 201 -842 0 FreeSans 160 0 0 0 M9
flabel metal2 917 -760 946 -738 0 FreeSans 160 0 0 0 D9
port 6 nsew
flabel metal1 698 -429 727 -361 0 FreeSans 160 0 0 0 GND
port 2 nsew
flabel metal1 918 -664 934 -657 0 FreeSans 160 0 0 0 D8
port 7 nsew
<< end >>
