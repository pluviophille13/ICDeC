magic
tech sky130A
timestamp 1729223146
<< nmos >>
rect -50 -40 50 40
<< ndiff >>
rect -79 34 -50 40
rect -79 -34 -73 34
rect -56 -34 -50 34
rect -79 -40 -50 -34
rect 50 34 79 40
rect 50 -34 56 34
rect 73 -34 79 34
rect 50 -40 79 -34
<< ndiffc >>
rect -73 -34 -56 34
rect 56 -34 73 34
<< poly >>
rect -50 76 50 84
rect -50 59 -42 76
rect 42 59 50 76
rect -50 40 50 59
rect -50 -59 50 -40
rect -50 -76 -42 -59
rect 42 -76 50 -59
rect -50 -84 50 -76
<< polycont >>
rect -42 59 42 76
rect -42 -76 42 -59
<< locali >>
rect -50 59 -42 76
rect 42 59 50 76
rect -73 34 -56 42
rect -73 -42 -56 -34
rect 56 34 73 42
rect 56 -42 73 -34
rect -50 -76 -42 -59
rect 42 -76 50 -59
<< viali >>
rect -42 59 42 76
rect -73 -34 -56 34
rect 56 -34 73 34
rect -42 -76 42 -59
<< metal1 >>
rect -48 76 48 79
rect -48 59 -42 76
rect 42 59 48 76
rect -48 56 48 59
rect -76 34 -53 40
rect -76 -34 -73 34
rect -56 -34 -53 34
rect -76 -40 -53 -34
rect 53 34 76 40
rect 53 -34 56 34
rect 73 -34 76 34
rect 53 -40 76 -34
rect -48 -59 48 -56
rect -48 -76 -42 -59
rect 42 -76 48 -59
rect -48 -79 48 -76
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.8 l 1 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 1 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
