magic
tech sky130A
magscale 1 2
timestamp 1729238107
<< nwell >>
rect -197 -1743 621 693
<< nsubdiff >>
rect -161 623 -101 657
rect 525 623 585 657
rect -161 597 -127 623
rect 551 597 585 623
rect -161 -1673 -127 -1647
rect 551 -1673 585 -1647
rect -161 -1707 -101 -1673
rect 525 -1707 585 -1673
<< nsubdiffcont >>
rect -101 623 525 657
rect -161 -1647 -127 597
rect 551 -1647 585 597
rect -101 -1707 525 -1673
<< poly >>
rect -6 52 24 57
rect -72 36 24 52
rect -72 2 -56 36
rect -22 2 24 36
rect -72 -14 24 2
rect 398 52 428 57
rect 398 36 494 52
rect 398 2 444 36
rect 478 2 494 36
rect 398 -14 494 2
rect -6 -413 24 -408
rect -72 -429 24 -413
rect -72 -463 -56 -429
rect -22 -463 24 -429
rect -72 -479 24 -463
rect 398 -413 428 -408
rect 398 -429 494 -413
rect 398 -463 444 -429
rect 478 -463 494 -429
rect -72 -561 24 -545
rect 82 -546 182 -478
rect 240 -546 340 -478
rect 398 -479 494 -463
rect -72 -595 -56 -561
rect -22 -595 24 -561
rect -72 -611 24 -595
rect -6 -616 24 -611
rect 398 -561 494 -545
rect 398 -595 444 -561
rect 478 -595 494 -561
rect 398 -611 494 -595
rect 398 -616 428 -611
rect -72 -1026 24 -1010
rect -72 -1060 -56 -1026
rect -22 -1060 24 -1026
rect -72 -1076 24 -1060
rect -6 -1081 24 -1076
rect 398 -1026 494 -1010
rect 398 -1060 444 -1026
rect 478 -1060 494 -1026
rect 398 -1076 494 -1060
rect 398 -1081 428 -1076
<< polycont >>
rect -56 2 -22 36
rect 444 2 478 36
rect -56 -463 -22 -429
rect 444 -463 478 -429
rect -56 -595 -22 -561
rect 444 -595 478 -561
rect -56 -1060 -22 -1026
rect 444 -1060 478 -1026
<< locali >>
rect -161 623 -101 657
rect 525 623 585 657
rect -161 597 -127 623
rect 551 597 585 623
rect -52 36 -18 83
rect 440 36 474 83
rect -72 2 -56 36
rect -22 2 -6 36
rect 428 2 444 36
rect 478 2 494 36
rect -52 -429 -18 -382
rect 440 -429 474 -382
rect -72 -463 -56 -429
rect -22 -463 -6 -429
rect 428 -463 444 -429
rect 478 -463 494 -429
rect -72 -595 -56 -561
rect -22 -595 -6 -561
rect 428 -595 444 -561
rect 478 -595 494 -561
rect -52 -642 -18 -595
rect 440 -642 474 -595
rect -72 -1060 -56 -1026
rect -22 -1060 -6 -1026
rect 428 -1060 444 -1026
rect 478 -1060 494 -1026
rect -52 -1107 -18 -1060
rect 440 -1107 474 -1060
rect -161 -1673 -127 -1647
rect 551 -1673 585 -1647
rect -161 -1707 -101 -1673
rect 525 -1707 585 -1673
<< viali >>
rect 150 623 268 657
rect -56 2 -22 36
rect 444 2 478 36
rect -56 -463 -22 -429
rect 444 -463 478 -429
rect -56 -595 -22 -561
rect 444 -595 478 -561
rect -56 -1060 -22 -1026
rect 444 -1060 478 -1026
<< metal1 >>
rect 138 657 280 663
rect 138 623 150 657
rect 268 623 280 657
rect 138 617 280 623
rect 429 588 489 594
rect -21 528 429 588
rect -21 95 39 528
rect 429 522 489 528
rect 175 95 185 271
rect 237 95 247 271
rect 377 95 387 271
rect 439 95 449 271
rect -58 42 -12 95
rect -68 36 -10 42
rect -68 2 -56 36
rect -22 2 -10 36
rect -68 -4 -10 2
rect 98 -35 166 2
rect 246 -7 256 45
rect 324 -7 334 45
rect 434 42 480 95
rect 432 36 490 42
rect 432 2 444 36
rect 478 2 490 36
rect 432 -4 490 2
rect 98 -64 324 -35
rect 88 -144 98 -92
rect 166 -144 176 -92
rect 256 -101 324 -64
rect -71 -370 -61 -194
rect -9 -370 70 -194
rect 175 -370 185 -194
rect 237 -370 247 -194
rect 352 -370 430 -194
rect 484 -370 494 -194
rect -58 -423 -12 -370
rect 434 -423 480 -370
rect -68 -429 -10 -423
rect -68 -463 -56 -429
rect -22 -463 -10 -429
rect -68 -469 -10 -463
rect 432 -429 490 -423
rect 432 -463 444 -429
rect 478 -463 490 -429
rect 432 -469 490 -463
rect -68 -561 -10 -555
rect -68 -595 -56 -561
rect -22 -595 -10 -561
rect -68 -601 -10 -595
rect 432 -561 490 -555
rect 432 -595 444 -561
rect 478 -595 490 -561
rect 432 -601 490 -595
rect -58 -654 -12 -601
rect 434 -654 480 -601
rect -71 -830 -61 -654
rect -9 -830 70 -654
rect 175 -830 185 -654
rect 237 -830 247 -654
rect 352 -830 430 -654
rect 484 -830 494 -654
rect 88 -932 98 -880
rect 166 -932 176 -880
rect 256 -960 324 -923
rect 98 -989 324 -960
rect -68 -1026 -10 -1020
rect 98 -1026 166 -989
rect -68 -1060 -56 -1026
rect -22 -1060 -10 -1026
rect -68 -1066 -10 -1060
rect -58 -1110 -12 -1066
rect 246 -1069 256 -1017
rect 324 -1069 334 -1017
rect 432 -1026 490 -1020
rect 432 -1060 444 -1026
rect 478 -1060 490 -1026
rect 432 -1066 490 -1060
rect 434 -1111 480 -1066
rect -52 -1295 70 -1119
rect 175 -1295 185 -1119
rect 237 -1295 247 -1119
rect 377 -1295 387 -1119
rect 439 -1295 449 -1119
rect -20 -1552 40 -1295
rect 429 -1552 489 -1546
rect -20 -1612 429 -1552
rect 429 -1618 489 -1612
<< via1 >>
rect 429 528 489 588
rect 185 95 237 271
rect 387 95 439 271
rect 256 -7 324 45
rect 98 -144 166 -92
rect -61 -370 -9 -194
rect 185 -370 237 -194
rect 430 -370 484 -194
rect -61 -830 -9 -654
rect 185 -830 237 -654
rect 430 -830 484 -654
rect 98 -932 166 -880
rect 256 -1069 324 -1017
rect 185 -1295 237 -1119
rect 387 -1295 439 -1119
rect 429 -1612 489 -1552
<< metal2 >>
rect 423 586 429 588
rect 489 586 495 588
rect 422 530 429 586
rect 489 530 496 586
rect 423 528 429 530
rect 489 528 495 530
rect -61 430 439 482
rect -61 -194 -9 430
rect 183 271 239 283
rect 183 86 239 95
rect 387 271 439 430
rect 185 85 237 86
rect 387 80 439 95
rect 256 45 324 51
rect 256 -37 324 -7
rect 98 -67 324 -37
rect 98 -92 166 -67
rect 98 -154 166 -144
rect -61 -654 -9 -370
rect 183 -194 239 -184
rect 183 -380 239 -370
rect 429 -194 485 -184
rect 429 -380 485 -370
rect -61 -1454 -9 -830
rect 183 -654 239 -644
rect 183 -840 239 -830
rect 429 -654 485 -644
rect 429 -840 485 -830
rect 98 -880 166 -870
rect 98 -957 166 -932
rect 98 -987 324 -957
rect 256 -1017 324 -987
rect 256 -1079 324 -1069
rect 183 -1119 239 -1104
rect 183 -1304 239 -1295
rect 387 -1119 439 -1104
rect 185 -1305 237 -1304
rect 387 -1454 439 -1295
rect -62 -1506 439 -1454
rect 423 -1554 429 -1552
rect 489 -1554 495 -1552
rect 422 -1610 429 -1554
rect 489 -1610 496 -1554
rect 423 -1612 429 -1610
rect 489 -1612 495 -1610
<< via2 >>
rect 431 530 487 586
rect 183 95 185 271
rect 185 95 237 271
rect 237 95 239 271
rect 183 -370 185 -194
rect 185 -370 237 -194
rect 237 -370 239 -194
rect 429 -370 430 -194
rect 430 -370 484 -194
rect 484 -370 485 -194
rect 183 -830 185 -654
rect 185 -830 237 -654
rect 237 -830 239 -654
rect 429 -830 430 -654
rect 430 -830 484 -654
rect 484 -830 485 -654
rect 183 -1295 185 -1119
rect 185 -1295 237 -1119
rect 237 -1295 239 -1119
rect 431 -1610 487 -1554
<< metal3 >>
rect 426 586 492 591
rect 426 530 431 586
rect 487 530 492 586
rect 426 525 492 530
rect 173 271 249 280
rect 173 95 183 271
rect 239 95 249 271
rect 173 -194 249 95
rect 429 -189 489 525
rect 173 -370 183 -194
rect 239 -370 249 -194
rect 173 -654 249 -370
rect 419 -194 495 -189
rect 419 -370 429 -194
rect 485 -370 495 -194
rect 419 -375 495 -370
rect 429 -649 489 -375
rect 173 -830 183 -654
rect 239 -830 249 -654
rect 173 -1119 249 -830
rect 419 -654 495 -649
rect 419 -830 429 -654
rect 485 -830 495 -654
rect 419 -835 495 -830
rect 173 -1295 183 -1119
rect 239 -1295 249 -1119
rect 173 -1304 249 -1295
rect 429 -1549 489 -835
rect 426 -1554 492 -1549
rect 426 -1610 431 -1554
rect 487 -1610 492 -1554
rect 426 -1615 492 -1610
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_0
timestamp 1729223943
transform 1 0 9 0 1 183
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_1
timestamp 1729223943
transform 1 0 413 0 1 183
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_2
timestamp 1729223943
transform 1 0 9 0 1 -1207
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_3
timestamp 1729223943
transform 1 0 9 0 1 -282
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_4
timestamp 1729223943
transform 1 0 413 0 1 -282
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_5
timestamp 1729223943
transform 1 0 413 0 1 -742
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_6
timestamp 1729223943
transform 1 0 413 0 1 -1207
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_7
timestamp 1729223943
transform 1 0 9 0 1 -742
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_BHVYY6  sky130_fd_pr__pfet_01v8_BHVYY6_0
timestamp 1729223943
transform 1 0 211 0 1 -1207
box -223 -200 223 200
use sky130_fd_pr__pfet_01v8_BHVYY6  sky130_fd_pr__pfet_01v8_BHVYY6_1
timestamp 1729223943
transform 1 0 211 0 1 183
box -223 -200 223 200
use sky130_fd_pr__pfet_01v8_BHVYY6  sky130_fd_pr__pfet_01v8_BHVYY6_2
timestamp 1729223943
transform 1 0 211 0 1 -282
box -223 -200 223 200
use sky130_fd_pr__pfet_01v8_BHVYY6  sky130_fd_pr__pfet_01v8_BHVYY6_3
timestamp 1729223943
transform 1 0 211 0 1 -742
box -223 -200 223 200
<< labels >>
flabel viali 206 640 206 640 0 FreeSans 1600 0 0 0 VDD
port 0 nsew
flabel metal3 461 497 461 497 0 FreeSans 1600 0 0 0 OUT
port 1 nsew
flabel metal2 80 454 80 454 0 FreeSans 1600 0 0 0 D6
port 2 nsew
flabel metal1 130 -27 130 -27 0 FreeSans 1600 0 0 0 VIP
port 3 nsew
flabel metal2 114 -76 114 -76 0 FreeSans 1600 0 0 0 VIN
port 4 nsew
flabel metal3 208 -508 208 -508 0 FreeSans 1600 0 0 0 D5
port 5 nsew
<< end >>
