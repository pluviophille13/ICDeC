magic
tech sky130A
timestamp 1729223146
<< nmos >>
rect -40 -50 40 50
<< ndiff >>
rect -69 44 -40 50
rect -69 -44 -63 44
rect -46 -44 -40 44
rect -69 -50 -40 -44
rect 40 44 69 50
rect 40 -44 46 44
rect 63 -44 69 44
rect 40 -50 69 -44
<< ndiffc >>
rect -63 -44 -46 44
rect 46 -44 63 44
<< poly >>
rect -40 86 40 94
rect -40 69 -32 86
rect 32 69 40 86
rect -40 50 40 69
rect -40 -69 40 -50
rect -40 -86 -32 -69
rect 32 -86 40 -69
rect -40 -94 40 -86
<< polycont >>
rect -32 69 32 86
rect -32 -86 32 -69
<< locali >>
rect -40 69 -32 86
rect 32 69 40 86
rect -63 44 -46 52
rect -63 -52 -46 -44
rect 46 44 63 52
rect 46 -52 63 -44
rect -40 -86 -32 -69
rect 32 -86 40 -69
<< viali >>
rect -32 69 32 86
rect -63 -44 -46 44
rect 46 -44 63 44
rect -32 -86 32 -69
<< metal1 >>
rect -38 86 38 89
rect -38 69 -32 86
rect 32 69 38 86
rect -38 66 38 69
rect -66 44 -43 50
rect -66 -44 -63 44
rect -46 -44 -43 44
rect -66 -50 -43 -44
rect 43 44 66 50
rect 43 -44 46 44
rect 63 -44 66 44
rect 43 -50 66 -44
rect -38 -69 38 -66
rect -38 -86 -32 -69
rect 32 -86 38 -69
rect -38 -89 38 -86
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1 l 0.8 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 1 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
